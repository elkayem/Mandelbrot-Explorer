
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_wild is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_wild;

architecture arch of colormap_wild is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"333",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed2",
      x"ed2",
      x"ed2",
      x"ed2",
      x"c57",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ed3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"ec3",
      x"eb3",
      x"eb3",
      x"eb4",
      x"eb4",
      x"eb4",
      x"eb4",
      x"eb4",
      x"eb4",
      x"eb4",
      x"eb4",
      x"db4",
      x"db4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da4",
      x"da5",
      x"da5",
      x"da5",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d95",
      x"d85",
      x"d85",
      x"d85",
      x"d85",
      x"d85",
      x"d86",
      x"d86",
      x"d86",
      x"d86",
      x"d86",
      x"d86",
      x"d86",
      x"c86",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c76",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c67",
      x"c57",
      x"c57",
      x"c57",
      x"10e",
      x"20e",
      x"20d",
      x"20d",
      x"20d",
      x"30d",
      x"30d",
      x"31d",
      x"31d",
      x"41c",
      x"41c",
      x"41c",
      x"41c",
      x"41c",
      x"51c",
      x"52c",
      x"52b",
      x"52b",
      x"62b",
      x"62b",
      x"62b",
      x"62b",
      x"62b",
      x"73a",
      x"73a",
      x"73a",
      x"73a",
      x"83a",
      x"83a",
      x"83a",
      x"839",
      x"849",
      x"949",
      x"949",
      x"949",
      x"949",
      x"a49",
      x"a48",
      x"a48",
      x"a58",
      x"a58",
      x"b58",
      x"b58",
      x"b58",
      x"b57",
      x"c57",
      x"c57",
      x"2d7",
      x"2d7",
      x"2d7",
      x"2d7",
      x"3d7",
      x"3c7",
      x"3c7",
      x"3c7",
      x"3c7",
      x"3c7",
      x"3c7",
      x"4c7",
      x"4c7",
      x"4c7",
      x"4b7",
      x"4b7",
      x"4b7",
      x"4b7",
      x"4b7",
      x"5b7",
      x"5b7",
      x"5b7",
      x"5b7",
      x"5b7",
      x"5a7",
      x"5a7",
      x"6a7",
      x"6a7",
      x"6a7",
      x"6a7",
      x"6a7",
      x"6a7",
      x"6a7",
      x"797",
      x"797",
      x"797",
      x"797",
      x"797",
      x"797",
      x"797",
      x"897",
      x"897",
      x"887",
      x"887",
      x"887",
      x"887",
      x"887",
      x"987",
      x"987",
      x"987",
      x"987",
      x"987",
      x"977",
      x"977",
      x"977",
      x"a77",
      x"a77",
      x"a77",
      x"a77",
      x"a77",
      x"a77",
      x"a67",
      x"b67",
      x"b67",
      x"b67",
      x"b67",
      x"b67",
      x"b67",
      x"b67",
      x"c67",
      x"c57",
      x"c57",
      x"e26",
      x"e26",
      x"e26",
      x"e26",
      x"e26",
      x"e26",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d46",
      x"d46",
      x"d46",
      x"d47",
      x"d47",
      x"d47",
      x"d47",
      x"d47",
      x"c47",
      x"c47"
   );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;