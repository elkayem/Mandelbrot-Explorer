
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_roygold is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_roygold;

architecture arch of colormap_roygold is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
     x"000",
      x"b69",
      x"b69",
      x"b69",
      x"b59",
      x"b59",
      x"b59",
      x"b59",
      x"b59",
      x"b58",
      x"b58",
      x"b58",
      x"b58",
      x"b48",
      x"a48",
      x"a48",
      x"a48",
      x"a48",
      x"a47",
      x"a47",
      x"a47",
      x"a37",
      x"a37",
      x"a37",
      x"a37",
      x"a37",
      x"a37",
      x"a36",
      x"a36",
      x"a36",
      x"a26",
      x"a26",
      x"a26",
      x"a26",
      x"a26",
      x"a26",
      x"a25",
      x"925",
      x"915",
      x"915",
      x"915",
      x"915",
      x"915",
      x"925",
      x"926",
      x"836",
      x"837",
      x"847",
      x"847",
      x"758",
      x"758",
      x"768",
      x"769",
      x"679",
      x"67a",
      x"68a",
      x"59a",
      x"59b",
      x"5ab",
      x"5ac",
      x"4bc",
      x"4bc",
      x"4cd",
      x"4cd",
      x"3de",
      x"3de",
      x"3ee",
      x"3ef",
      x"2ff",
      x"2ff",
      x"2ff",
      x"2ff",
      x"2ee",
      x"2ee",
      x"2ee",
      x"2ed",
      x"2dd",
      x"2dd",
      x"2dc",
      x"2dc",
      x"2cc",
      x"2cb",
      x"2cb",
      x"2cb",
      x"2ca",
      x"2ba",
      x"2ba",
      x"1b9",
      x"1b9",
      x"1a9",
      x"1a8",
      x"1a8",
      x"1a8",
      x"197",
      x"197",
      x"197",
      x"196",
      x"186",
      x"186",
      x"185",
      x"185",
      x"185",
      x"174",
      x"174",
      x"174",
      x"173",
      x"163",
      x"163",
      x"162",
      x"162",
      x"152",
      x"151",
      x"151",
      x"151",
      x"151",
      x"151",
      x"151",
      x"152",
      x"142",
      x"142",
      x"242",
      x"242",
      x"242",
      x"242",
      x"242",
      x"243",
      x"243",
      x"243",
      x"243",
      x"243",
      x"243",
      x"243",
      x"244",
      x"344",
      x"334",
      x"334",
      x"334",
      x"334",
      x"334",
      x"335",
      x"335",
      x"335",
      x"335",
      x"335",
      x"335",
      x"335",
      x"335",
      x"435",
      x"435",
      x"545",
      x"545",
      x"645",
      x"644",
      x"654",
      x"754",
      x"754",
      x"854",
      x"864",
      x"963",
      x"963",
      x"963",
      x"a73",
      x"a73",
      x"b73",
      x"b73",
      x"c82",
      x"c82",
      x"c82",
      x"d82",
      x"d92",
      x"e92",
      x"e92",
      x"f91",
      x"f91",
      x"f91",
      x"e91",
      x"e91",
      x"e91",
      x"e81",
      x"d81",
      x"d81",
      x"d81",
      x"d81",
      x"c81",
      x"c71",
      x"c71",
      x"c71",
      x"b71",
      x"b71",
      x"b71",
      x"b61",
      x"a61",
      x"a61",
      x"a61",
      x"a61",
      x"961",
      x"961",
      x"951",
      x"950",
      x"850",
      x"850",
      x"850",
      x"850",
      x"740",
      x"740",
      x"740",
      x"740",
      x"640",
      x"640",
      x"630",
      x"630",
      x"530",
      x"530",
      x"530",
      x"630",
      x"631",
      x"641",
      x"741",
      x"741",
      x"842",
      x"852",
      x"852",
      x"952",
      x"953",
      x"a53",
      x"a63",
      x"b63",
      x"b64",
      x"b64",
      x"c64",
      x"c74",
      x"d75",
      x"d75",
      x"d75",
      x"e85",
      x"e86",
      x"f86",
      x"f86",
      x"e86",
      x"e86",
      x"e87",
      x"d87",
      x"d97",
      x"c97",
      x"c98",
      x"c98",
      x"b98",
      x"b98",
      x"a99",
      x"a99",
      x"999",
      x"999",
      x"99a",
      x"89a",
      x"89a",
      x"79a"
   );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;