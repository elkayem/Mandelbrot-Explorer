
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_polar is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_polar;

architecture arch of colormap_polar is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"000",
      x"ead",
      x"ead",
      x"ead",
      x"ead",
      x"ebc",
      x"ebc",
      x"ebc",
      x"ebb",
      x"ecb",
      x"ecb",
      x"ecb",
      x"dda",
      x"cda",
      x"ada",
      x"8da",
      x"7ea",
      x"5ea",
      x"3ea",
      x"4ea",
      x"4ea",
      x"5da",
      x"5da",
      x"6da",
      x"6db",
      x"6cb",
      x"7cb",
      x"7cb",
      x"8cb",
      x"8bb",
      x"9bc",
      x"6d8",
      x"0ee",
      x"1ee",
      x"1de",
      x"1de",
      x"1de",
      x"2de",
      x"2cd",
      x"2cd",
      x"2cd",
      x"3bd",
      x"3bd",
      x"3bd",
      x"3bc",
      x"4ac",
      x"4ac",
      x"4ac",
      x"49c",
      x"59c",
      x"59c",
      x"59b",
      x"58b",
      x"68b",
      x"68b",
      x"68b",
      x"68b",
      x"78b",
      x"79b",
      x"79b",
      x"79a",
      x"8aa",
      x"8aa",
      x"8aa",
      x"8aa",
      x"9ba",
      x"9ba",
      x"9ba",
      x"9ca",
      x"aca",
      x"aca",
      x"aca",
      x"bd9",
      x"bd9",
      x"bc9",
      x"bc9",
      x"bc9",
      x"bc9",
      x"bb9",
      x"bb9",
      x"bb9",
      x"bb9",
      x"baa",
      x"baa",
      x"caa",
      x"c9a",
      x"c9a",
      x"c9a",
      x"c9a",
      x"c8a",
      x"c8a",
      x"c8a",
      x"c7a",
      x"c7a",
      x"c8a",
      x"c89",
      x"d89",
      x"d89",
      x"d89",
      x"d89",
      x"d89",
      x"d88",
      x"d98",
      x"d98",
      x"d98",
      x"d98",
      x"d97",
      x"d97",
      x"d97",
      x"e97",
      x"ea7",
      x"ea6",
      x"ea6",
      x"ea6",
      x"ea6",
      x"ea6",
      x"da6",
      x"ca7",
      x"ba7",
      x"a98",
      x"a98",
      x"999",
      x"89a",
      x"78a",
      x"899",
      x"9a7",
      x"bb5",
      x"cc3",
      x"ed1",
      x"dc1",
      x"dc1",
      x"cb1",
      x"ca1",
      x"ca1",
      x"b91",
      x"b81",
      x"a71",
      x"a71",
      x"961",
      x"951",
      x"951",
      x"841",
      x"831",
      x"731",
      x"721",
      x"611",
      x"622",
      x"623",
      x"533",
      x"534",
      x"445",
      x"456",
      x"357",
      x"368",
      x"269",
      x"27a",
      x"28a",
      x"18b",
      x"19c",
      x"0ad",
      x"19d",
      x"29d",
      x"28d",
      x"38d",
      x"47e",
      x"57e",
      x"56e",
      x"66e",
      x"75e",
      x"85e",
      x"85e",
      x"94e",
      x"a4e",
      x"b3e",
      x"b3f",
      x"c2f",
      x"d2f",
      x"e1f",
      x"f1f",
      x"e1f",
      x"d1f",
      x"c1e",
      x"b1e",
      x"91e",
      x"81e",
      x"72d",
      x"62d",
      x"52d",
      x"42d",
      x"32c",
      x"22c",
      x"13c",
      x"23c",
      x"24c",
      x"35b",
      x"45b",
      x"56b",
      x"67b",
      x"68b",
      x"78a",
      x"89a",
      x"9aa",
      x"999",
      x"999",
      x"988",
      x"987",
      x"a76",
      x"a76",
      x"a65",
      x"a64",
      x"a53",
      x"a53",
      x"a42",
      x"b41",
      x"b30",
      x"b31",
      x"a32",
      x"a42",
      x"a43",
      x"943",
      x"944",
      x"945",
      x"845",
      x"846",
      x"847",
      x"747",
      x"758",
      x"758",
      x"659",
      x"659",
      x"759",
      x"75a",
      x"85a",
      x"85a",
      x"85a",
      x"95a",
      x"94b",
      x"94b",
      x"a4b",
      x"a4b",
      x"b4b",
      x"b4c",
      x"b4c",
      x"c4c",
      x"c4c",
      x"d4c",
      x"d4c",
      x"d4d",
      x"e4d",
      x"e4d",
      x"f3d",
      x"e3d",
      x"e3d",
      x"e3c",
      x"e3c",
      x"d3b"
   );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;