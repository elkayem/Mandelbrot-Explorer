
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_caramel is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_caramel;

architecture arch of colormap_caramel is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"333",
      x"a8c",
      x"a8c",
      x"b9c",
      x"b9c",
      x"c9c",
      x"c9c",
      x"d9c",
      x"dac",
      x"eac",
      x"eac",
      x"eab",
      x"d9b",
      x"c8b",
      x"c7b",
      x"b7a",
      x"a6a",
      x"95a",
      x"959",
      x"849",
      x"739",
      x"858",
      x"a78",
      x"b98",
      x"cb7",
      x"ed7",
      x"dc7",
      x"cb8",
      x"bb9",
      x"aa9",
      x"99a",
      x"89b",
      x"88b",
      x"77c",
      x"67d",
      x"67c",
      x"77a",
      x"879",
      x"978",
      x"a76",
      x"b75",
      x"c74",
      x"d82",
      x"d82",
      x"d83",
      x"d83",
      x"d83",
      x"d93",
      x"d94",
      x"d94",
      x"d94",
      x"d94",
      x"da5",
      x"da5",
      x"da5",
      x"ea5",
      x"ea6",
      x"eb6",
      x"eb6",
      x"eb6",
      x"eb7",
      x"eb7",
      x"ec7",
      x"ec7",
      x"ec8",
      x"ec8",
      x"ed8",
      x"ed8",
      x"ed8",
      x"ec8",
      x"dc8",
      x"dc8",
      x"cb8",
      x"cb8",
      x"bb8",
      x"ba8",
      x"aa8",
      x"aa8",
      x"998",
      x"998",
      x"997",
      x"887",
      x"887",
      x"787",
      x"777",
      x"677",
      x"677",
      x"567",
      x"567",
      x"467",
      x"457",
      x"357",
      x"346",
      x"356",
      x"356",
      x"466",
      x"466",
      x"466",
      x"576",
      x"576",
      x"586",
      x"686",
      x"696",
      x"696",
      x"796",
      x"7a6",
      x"7a6",
      x"8b6",
      x"8b6",
      x"8b6",
      x"9c6",
      x"9c6",
      x"9d6",
      x"9d6",
      x"9c6",
      x"9c6",
      x"9c6",
      x"9c5",
      x"9b5",
      x"9b5",
      x"9b5",
      x"9b5",
      x"9a5",
      x"9a5",
      x"9a5",
      x"9a4",
      x"994",
      x"994",
      x"994",
      x"994",
      x"984",
      x"984",
      x"984",
      x"973",
      x"a74",
      x"a85",
      x"a86",
      x"b87",
      x"b87",
      x"b88",
      x"b99",
      x"c9a",
      x"c9a",
      x"c9a",
      x"c99",
      x"c99",
      x"c89",
      x"c89",
      x"c88",
      x"c88",
      x"c88",
      x"b88",
      x"b87",
      x"b87",
      x"b87",
      x"b87",
      x"b76",
      x"b76",
      x"b76",
      x"b76",
      x"b76",
      x"b75",
      x"b75",
      x"b75",
      x"b75",
      x"b74",
      x"b64",
      x"b64",
      x"b64",
      x"a63",
      x"a63",
      x"a63",
      x"a63",
      x"a62",
      x"a62",
      x"963",
      x"863",
      x"863",
      x"763",
      x"763",
      x"664",
      x"564",
      x"564",
      x"464",
      x"365",
      x"375",
      x"275",
      x"275",
      x"175",
      x"076",
      x"076",
      x"076",
      x"076",
      x"076",
      x"076",
      x"066",
      x"066",
      x"066",
      x"067",
      x"067",
      x"067",
      x"057",
      x"057",
      x"057",
      x"057",
      x"057",
      x"047",
      x"047",
      x"048",
      x"048",
      x"048",
      x"048",
      x"038",
      x"038",
      x"138",
      x"348",
      x"449",
      x"559",
      x"759",
      x"869",
      x"a6a",
      x"b6a",
      x"c7a",
      x"c7a",
      x"c7a",
      x"c7a",
      x"c8a",
      x"c8a",
      x"c8a",
      x"c8a",
      x"c8a",
      x"c8a",
      x"c9a",
      x"b9a",
      x"b9a",
      x"b9a",
      x"b9a",
      x"baa",
      x"baa",
      x"baa",
      x"baa",
      x"baa",
      x"bba",
      x"aba",
      x"aba",
      x"aba",
      x"aba",
      x"aca",
      x"aca",
      x"aca",
      x"aca",
      x"aca",
      x"ada",
      x"9da",
      x"9da",
      x"8db"
   );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;