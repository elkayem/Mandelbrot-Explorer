
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_tropic is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_tropic;

architecture arch of colormap_tropic is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"000",
      x"fbc",
      x"ebc",
      x"dbc",
      x"dbb",
      x"cbb",
      x"bbb",
      x"bbb",
      x"aab",
      x"9aa",
      x"9aa",
      x"8aa",
      x"7aa",
      x"7aa",
      x"7a9",
      x"7a9",
      x"7a9",
      x"7a9",
      x"7a9",
      x"8a9",
      x"8a9",
      x"8a9",
      x"8a9",
      x"8a9",
      x"8a9",
      x"999",
      x"999",
      x"999",
      x"999",
      x"999",
      x"999",
      x"999",
      x"a99",
      x"a99",
      x"a99",
      x"a99",
      x"a9a",
      x"a9a",
      x"a9a",
      x"99a",
      x"99a",
      x"99a",
      x"99a",
      x"99a",
      x"99a",
      x"99a",
      x"99a",
      x"99b",
      x"99b",
      x"99b",
      x"99b",
      x"89b",
      x"89b",
      x"89b",
      x"89b",
      x"89b",
      x"89b",
      x"89b",
      x"89b",
      x"89c",
      x"89c",
      x"89c",
      x"89c",
      x"79c",
      x"79c",
      x"79c",
      x"79c",
      x"79c",
      x"79c",
      x"79c",
      x"79d",
      x"79d",
      x"79d",
      x"79d",
      x"79d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"69d",
      x"6ad",
      x"6ad",
      x"6ad",
      x"6ad",
      x"6ad",
      x"6ad",
      x"6ad",
      x"6ad",
      x"5bd",
      x"5bd",
      x"5bd",
      x"5bd",
      x"5bd",
      x"5bd",
      x"5bd",
      x"5cc",
      x"5cc",
      x"5cc",
      x"5cc",
      x"5cc",
      x"5cc",
      x"5cc",
      x"5cc",
      x"5dc",
      x"5dc",
      x"5dc",
      x"5dc",
      x"5dc",
      x"5dc",
      x"5dc",
      x"5ec",
      x"5ec",
      x"5ec",
      x"5ec",
      x"5ec",
      x"4ec",
      x"4ec",
      x"4ec",
      x"4fc",
      x"4fc",
      x"4fc",
      x"4fc",
      x"6fa",
      x"8e8",
      x"ae6",
      x"ce4",
      x"ee2",
      x"ed2",
      x"dd3",
      x"dd4",
      x"dd4",
      x"dc5",
      x"dc6",
      x"cc6",
      x"cc7",
      x"cb8",
      x"cb8",
      x"cb9",
      x"bb9",
      x"baa",
      x"bab",
      x"bab",
      x"bac",
      x"998",
      x"885",
      x"772",
      x"772",
      x"763",
      x"863",
      x"863",
      x"863",
      x"854",
      x"854",
      x"854",
      x"955",
      x"945",
      x"945",
      x"945",
      x"946",
      x"936",
      x"a36",
      x"a37",
      x"a37",
      x"a27",
      x"a27",
      x"a28",
      x"a27",
      x"a37",
      x"937",
      x"937",
      x"947",
      x"947",
      x"847",
      x"857",
      x"857",
      x"857",
      x"767",
      x"767",
      x"767",
      x"777",
      x"677",
      x"677",
      x"687",
      x"587",
      x"587",
      x"597",
      x"597",
      x"497",
      x"4a7",
      x"4a7",
      x"4a7",
      x"3b7",
      x"3b7",
      x"3b7",
      x"3b7",
      x"3b7",
      x"4a7",
      x"4a7",
      x"4a7",
      x"4a7",
      x"597",
      x"597",
      x"597",
      x"597",
      x"596",
      x"686",
      x"686",
      x"686",
      x"686",
      x"676",
      x"776",
      x"776",
      x"776",
      x"776",
      x"866",
      x"866",
      x"866",
      x"866",
      x"855",
      x"955",
      x"955",
      x"955",
      x"955",
      x"945",
      x"a45",
      x"a45",
      x"a45",
      x"a35",
      x"b35",
      x"b35",
      x"b35",
      x"b35",
      x"b24",
      x"c24",
      x"c24",
      x"c24",
      x"c14",
      x"d14",
      x"d14",
      x"c24",
      x"c24",
      x"c24",
      x"c24",
      x"c34",
      x"c34",
      x"b35",
      x"b35",
      x"b45",
      x"b45"
	  );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;