
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_rose1 is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_rose1;

architecture arch of colormap_rose1 is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"000",
      x"7cd",
      x"7cd",
      x"7cd",
      x"7dd",
      x"8dd",
      x"8cc",
      x"8bc",
      x"8ab",
      x"89b",
      x"99b",
      x"98a",
      x"97a",
      x"969",
      x"a69",
      x"a58",
      x"a48",
      x"a38",
      x"b37",
      x"b27",
      x"a37",
      x"a36",
      x"935",
      x"935",
      x"934",
      x"834",
      x"833",
      x"732",
      x"732",
      x"731",
      x"631",
      x"630",
      x"732",
      x"732",
      x"732",
      x"722",
      x"722",
      x"722",
      x"722",
      x"622",
      x"622",
      x"622",
      x"621",
      x"621",
      x"621",
      x"621",
      x"621",
      x"621",
      x"621",
      x"621",
      x"611",
      x"611",
      x"611",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"511",
      x"500",
      x"500",
      x"500",
      x"500",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"400",
      x"500",
      x"501",
      x"501",
      x"501",
      x"501",
      x"501",
      x"501",
      x"601",
      x"601",
      x"602",
      x"602",
      x"602",
      x"602",
      x"602",
      x"602",
      x"702",
      x"702",
      x"703",
      x"703",
      x"703",
      x"703",
      x"703",
      x"803",
      x"803",
      x"803",
      x"804",
      x"804",
      x"804",
      x"804",
      x"904",
      x"904",
      x"904",
      x"904",
      x"904",
      x"905",
      x"905",
      x"905",
      x"a05",
      x"a05",
      x"a05",
      x"a05",
      x"a05",
      x"a06",
      x"a06",
      x"b06",
      x"b06",
      x"b06",
      x"b06",
      x"b06",
      x"b06",
      x"b07",
      x"c07",
      x"c07",
      x"c07",
      x"c07",
      x"c07",
      x"c07",
      x"c07",
      x"c08",
      x"d08",
      x"d08",
      x"d08",
      x"d18",
      x"d17",
      x"d17",
      x"d27",
      x"d27",
      x"d26",
      x"d36",
      x"d36",
      x"d46",
      x"d45",
      x"d55",
      x"d55",
      x"d55",
      x"d64",
      x"d64",
      x"d74",
      x"e73",
      x"e83",
      x"e83",
      x"e93",
      x"e92",
      x"e92",
      x"ea2",
      x"ea2",
      x"eb1",
      x"eb1",
      x"ec1",
      x"ec0",
      x"ec0",
      x"ec1",
      x"ec1",
      x"ec1",
      x"ec1",
      x"ec1",
      x"ec1",
      x"ec1",
      x"ec1",
      x"dc2",
      x"dc2",
      x"dc2",
      x"dc2",
      x"dc2",
      x"dc2",
      x"dc2",
      x"dc2",
      x"dc3",
      x"cb3",
      x"cb3",
      x"cb3",
      x"cb3",
      x"cb3",
      x"cb3",
      x"cb3",
      x"cb4",
      x"cb4",
      x"bb4",
      x"bb4",
      x"bb4",
      x"bb4",
      x"bb4",
      x"bb4",
      x"bb5",
      x"bb5",
      x"bb5",
      x"ab5",
      x"ab5",
      x"ab5",
      x"ab5",
      x"ab5",
      x"ab6",
      x"ab6",
      x"aa6",
      x"aa6",
      x"9a6",
      x"9a6",
      x"9a6",
      x"9a6",
      x"9a7",
      x"9a7",
      x"9a7",
      x"9a7",
      x"9a7",
      x"8a7",
      x"8a7",
      x"8a7",
      x"8a8",
      x"8a8",
      x"8a8",
      x"8a8",
      x"8a8",
      x"8a8",
      x"7a8",
      x"7a8",
      x"7a9",
      x"7a9",
      x"7a9",
      x"799",
      x"799",
      x"74d",
      x"75d",
      x"75d",
      x"75d",
      x"76d",
      x"76d",
      x"77d",
      x"77d",
      x"78d",
      x"78d",
      x"78d",
      x"79d",
      x"79d",
      x"7ad",
      x"7ad",
      x"7bd",
      x"7bd"
	  );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;