
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_candy is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_candy;

architecture arch of colormap_candy is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"000",
      x"c82",
      x"c92",
      x"c92",
      x"c92",
      x"d92",
      x"d92",
      x"d92",
      x"d92",
      x"da2",
      x"ea2",
      x"ea1",
      x"ea1",
      x"ea1",
      x"ea1",
      x"ea1",
      x"fa1",
      x"fb1",
      x"fb1",
      x"fb1",
      x"fb1",
      x"fb1",
      x"fa2",
      x"fa2",
      x"fa2",
      x"f92",
      x"f92",
      x"f92",
      x"f82",
      x"f83",
      x"f83",
      x"f73",
      x"f73",
      x"f73",
      x"f73",
      x"f64",
      x"f64",
      x"f64",
      x"f54",
      x"f54",
      x"f54",
      x"f45",
      x"f45",
      x"f45",
      x"f35",
      x"f35",
      x"f35",
      x"f25",
      x"f26",
      x"f26",
      x"e36",
      x"d46",
      x"c56",
      x"a66",
      x"987",
      x"897",
      x"7a7",
      x"6b7",
      x"5d7",
      x"f0f",
      x"e2d",
      x"c5c",
      x"a8b",
      x"9b9",
      x"7e8",
      x"9b9",
      x"9b9",
      x"9b9",
      x"ab8",
      x"ab8",
      x"ac8",
      x"bc7",
      x"bc7",
      x"bc7",
      x"cc6",
      x"cc6",
      x"cc6",
      x"dd6",
      x"dd5",
      x"dd5",
      x"ed5",
      x"ed4",
      x"ed4",
      x"fd4",
      x"fd3",
      x"fe3",
      x"fe3",
      x"fe3",
      x"fe2",
      x"fe3",
      x"fe3",
      x"fe3",
      x"fe3",
      x"fd3",
      x"fd3",
      x"fd3",
      x"fd3",
      x"fd3",
      x"fd3",
      x"fd4",
      x"fd4",
      x"fc4",
      x"fc4",
      x"fc4",
      x"fc4",
      x"ec4",
      x"ec4",
      x"ec4",
      x"ec4",
      x"eb5",
      x"eb5",
      x"eb5",
      x"eb5",
      x"eb5",
      x"eb5",
      x"eb5",
      x"db5",
      x"db5",
      x"da5",
      x"da5",
      x"da6",
      x"da6",
      x"da6",
      x"da6",
      x"da6",
      x"da6",
      x"c96",
      x"c96",
      x"c96",
      x"c96",
      x"c97",
      x"c97",
      x"c97",
      x"c97",
      x"c97",
      x"c87",
      x"c87",
      x"b87",
      x"b87",
      x"b87",
      x"b87",
      x"b88",
      x"b88",
      x"b78",
      x"b78",
      x"b78",
      x"b78",
      x"b78",
      x"a78",
      x"a78",
      x"a78",
      x"a69",
      x"a69",
      x"a69",
      x"a69",
      x"a69",
      x"a69",
      x"a69",
      x"a69",
      x"969",
      x"959",
      x"959",
      x"95a",
      x"95a",
      x"95a",
      x"95a",
      x"95a",
      x"95a",
      x"94a",
      x"94a",
      x"84a",
      x"84a",
      x"84b",
      x"84a",
      x"84a",
      x"83a",
      x"83a",
      x"82a",
      x"829",
      x"829",
      x"819",
      x"819",
      x"819",
      x"809",
      x"808",
      x"809",
      x"819",
      x"819",
      x"819",
      x"819",
      x"818",
      x"818",
      x"818",
      x"818",
      x"828",
      x"828",
      x"828",
      x"828",
      x"828",
      x"828",
      x"828",
      x"828",
      x"838",
      x"838",
      x"838",
      x"838",
      x"838",
      x"838",
      x"838",
      x"838",
      x"848",
      x"848",
      x"547",
      x"547",
      x"547",
      x"547",
      x"547",
      x"547",
      x"557",
      x"557",
      x"557",
      x"557",
      x"557",
      x"557",
      x"557",
      x"567",
      x"567",
      x"567",
      x"567",
      x"567",
      x"567",
      x"567",
      x"567",
      x"577",
      x"577",
      x"576",
      x"576",
      x"576",
      x"576",
      x"576",
      x"576",
      x"586",
      x"586",
      x"586",
      x"586",
      x"586",
      x"586",
      x"586",
      x"586",
      x"596",
      x"596",
      x"596",
      x"596",
      x"596",
      x"596",
      x"596"
	  );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;