
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_rosewht is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_rosewht;

architecture arch of colormap_rosewht is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"000",
      x"fc9",
      x"fc9",
      x"fc9",
      x"fc9",
      x"fc9",
      x"fc9",
      x"fc9",
      x"fc9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fd9",
      x"fe8",
      x"fe8",
      x"fe8",
      x"fe8",
      x"fe8",
      x"fe8",
      x"fe8",
      x"fe8",
      x"fe8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff8",
      x"ff9",
      x"ff9",
      x"ff9",
      x"ff9",
      x"ff9",
      x"ffa",
      x"ffa",
      x"ffa",
      x"ffa",
      x"ffb",
      x"ffb",
      x"ffb",
      x"ffb",
      x"ffb",
      x"ffc",
      x"ffc",
      x"ffc",
      x"ffc",
      x"ffc",
      x"ffd",
      x"ffd",
      x"ffd",
      x"ffd",
      x"ffe",
      x"ffe",
      x"ffe",
      x"ffe",
      x"ffe",
      x"fff",
      x"fff",
      x"fff",
      x"ffe",
      x"fee",
      x"fee",
      x"fed",
      x"fdd",
      x"fdd",
      x"fdc",
      x"ecc",
      x"ecc",
      x"ecb",
      x"dcb",
      x"dbb",
      x"dba",
      x"cba",
      x"caa",
      x"ca9",
      x"ba9",
      x"b99",
      x"b98",
      x"a98",
      x"a88",
      x"a87",
      x"987",
      x"977",
      x"876",
      x"866",
      x"766",
      x"655",
      x"655",
      x"545",
      x"444",
      x"445",
      x"545",
      x"545",
      x"535",
      x"535",
      x"635",
      x"635",
      x"735",
      x"735",
      x"835",
      x"835",
      x"825",
      x"835",
      x"835",
      x"835",
      x"945",
      x"945",
      x"945",
      x"945",
      x"955",
      x"955",
      x"945",
      x"945",
      x"a45",
      x"a45",
      x"a45",
      x"a45",
      x"a45",
      x"a45",
      x"a45",
      x"a45",
      x"a45",
      x"b45",
      x"b46",
      x"b46",
      x"b46",
      x"b46",
      x"b46",
      x"b46",
      x"b46",
      x"c46",
      x"c46",
      x"c46",
      x"c46",
      x"c46",
      x"c46",
      x"c46",
      x"c46",
      x"c46",
      x"d46",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"d36",
      x"e46",
      x"e46",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e47",
      x"e48",
      x"e48",
      x"e58",
      x"e58",
      x"e58",
      x"e58",
      x"e58",
      x"e58",
      x"e58",
      x"e58",
      x"e59",
      x"e59",
      x"e59",
      x"e59",
      x"e59",
      x"e59",
      x"e59",
      x"f59",
      x"f69",
      x"f69",
      x"f69",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6a",
      x"f6b",
      x"f6b",
      x"f7b",
      x"f7b",
      x"f7b",
      x"f7b",
      x"f7b",
      x"f7b",
      x"f7b",
      x"f7b",
      x"f7c",
      x"f7c",
      x"f7c",
      x"f7c",
      x"f7c",
      x"f7c",
      x"f7c",
      x"f8c",
      x"f8c",
      x"f8c",
      x"f8c",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8d",
      x"f8e",
      x"f8e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9e",
      x"f9f",
      x"f9f",
      x"f9f",
      x"f9f",
      x"f9f",
      x"f9f",
      x"f9f",
      x"faf",
      x"faf",
      x"faf"
	  );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;