
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity colormap_stargate is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(11 downto 0)
   );
end colormap_stargate;

architecture arch of colormap_stargate is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=12;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant colormap: rom_type:=(  -- 2^4-by-12
      x"000",
      x"69e",
      x"79e",
      x"79e",
      x"7ad",
      x"8ad",
      x"8ad",
      x"8ad",
      x"8bc",
      x"8bc",
      x"8bc",
      x"8bc",
      x"8bb",
      x"8bb",
      x"8cb",
      x"8cb",
      x"9ca",
      x"9ca",
      x"9ca",
      x"9ca",
      x"9ca",
      x"9ca",
      x"9da",
      x"9da",
      x"9da",
      x"9da",
      x"9da",
      x"9da",
      x"9ea",
      x"aea",
      x"aea",
      x"aea",
      x"aea",
      x"aea",
      x"aea",
      x"afa",
      x"afa",
      x"afa",
      x"afa",
      x"afa",
      x"afa",
      x"afa",
      x"afa",
      x"afa",
      x"bfa",
      x"bea",
      x"bea",
      x"bea",
      x"beb",
      x"bdb",
      x"adb",
      x"adb",
      x"adb",
      x"bcb",
      x"bcb",
      x"ccb",
      x"ccb",
      x"dbb",
      x"dbb",
      x"ebb",
      x"fbb",
      x"fbb",
      x"fbb",
      x"fab",
      x"fab",
      x"fab",
      x"fab",
      x"fab",
      x"fab",
      x"fab",
      x"eab",
      x"e9b",
      x"e9b",
      x"e9b",
      x"e9b",
      x"d9b",
      x"d9b",
      x"d9b",
      x"d9b",
      x"d8b",
      x"d8b",
      x"d8b",
      x"d8b",
      x"d8b",
      x"d8b",
      x"d8c",
      x"d8c",
      x"d7b",
      x"d7b",
      x"d7b",
      x"e7b",
      x"e7b",
      x"e7a",
      x"e7a",
      x"e7a",
      x"e6a",
      x"e69",
      x"e69",
      x"e69",
      x"e69",
      x"e58",
      x"e58",
      x"e58",
      x"e58",
      x"e49",
      x"e49",
      x"e59",
      x"e59",
      x"e6a",
      x"e6a",
      x"e7a",
      x"e7a",
      x"e8b",
      x"e8b",
      x"f9b",
      x"fab",
      x"fbc",
      x"fcc",
      x"fdc",
      x"feb",
      x"ffb",
      x"ffb",
      x"ffb",
      x"ffb",
      x"ffb",
      x"fea",
      x"fea",
      x"fea",
      x"fea",
      x"fda",
      x"fda",
      x"fda",
      x"fda",
      x"fca",
      x"fca",
      x"fca",
      x"fca",
      x"fca",
      x"fca",
      x"fca",
      x"fda",
      x"fda",
      x"fd9",
      x"fda",
      x"fda",
      x"fda",
      x"edb",
      x"edb",
      x"edb",
      x"edb",
      x"edb",
      x"edb",
      x"ecb",
      x"ecb",
      x"dcb",
      x"dcb",
      x"dcb",
      x"dcb",
      x"dcb",
      x"dcb",
      x"dcb",
      x"dba",
      x"cba",
      x"cba",
      x"cba",
      x"cba",
      x"cba",
      x"cba",
      x"cba",
      x"caa",
      x"baa",
      x"baa",
      x"baa",
      x"baa",
      x"baa",
      x"baa",
      x"b9a",
      x"b9a",
      x"b9a",
      x"a99",
      x"a99",
      x"a99",
      x"a99",
      x"a99",
      x"a89",
      x"a89",
      x"a89",
      x"989",
      x"989",
      x"989",
      x"989",
      x"989",
      x"989",
      x"979",
      x"979",
      x"879",
      x"879",
      x"878",
      x"878",
      x"878",
      x"868",
      x"868",
      x"868",
      x"768",
      x"768",
      x"768",
      x"768",
      x"767",
      x"767",
      x"767",
      x"667",
      x"656",
      x"656",
      x"656",
      x"656",
      x"655",
      x"656",
      x"656",
      x"556",
      x"556",
      x"556",
      x"546",
      x"547",
      x"547",
      x"547",
      x"547",
      x"448",
      x"448",
      x"448",
      x"448",
      x"349",
      x"349",
      x"359",
      x"35a",
      x"35a",
      x"35a",
      x"25a",
      x"25b",
      x"36b",
      x"36b",
      x"36b",
      x"36c",
      x"36c",
      x"37d",
      x"37d",
      x"37e",
      x"37e",
      x"47e",
      x"48e",
      x"48f",
      x"48f",
      x"58f",
      x"58f",
      x"69e",
      x"38e",
      x"38e"
	  );
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= colormap(to_integer(unsigned(addr_reg)));
end arch;